library IEEE;
use IEEE.numeric_std.all;

package custom_types is
    
    type integer_array is array (natural range <>) of integer;
    
end package custom_types;